/*
    Neptune v1.2.0 proportional window, for tinytapeout3.
    Copyright (C) 2023 Pat Deegan, https://psychogenic.com
    This program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.
    This program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.
    You should have received a copy of the GNU General Public License
    along with this program.  If not, see <https://www.gnu.org/licenses/>.
*/

`default_nettype none
`timescale 1ns/1ps
/* Generated by Yosys 0.28+1 (git sha1 a9c792dce, clang 10.0.0-4ubuntu1 -fPIC -Os) */

module discriminator(rst, clk, edge_count, note, match_high, match_far, match_exact);
  reg \$auto$verilog_backend.cc:2097:dump_module$5  = 0;
  wire \$1 ;
  wire [3:0] \$100 ;
  wire [3:0] \$102 ;
  wire [3:0] \$104 ;
  wire [3:0] \$106 ;
  wire [3:0] \$108 ;
  wire \$11 ;
  wire \$110 ;
  wire [8:0] \$112 ;
  wire \$114 ;
  wire [8:0] \$116 ;
  wire \$118 ;
  wire [8:0] \$120 ;
  wire \$122 ;
  wire [8:0] \$124 ;
  wire \$126 ;
  wire [8:0] \$128 ;
  wire \$13 ;
  wire \$130 ;
  wire [8:0] \$132 ;
  wire \$134 ;
  wire [8:0] \$136 ;
  wire \$138 ;
  wire [8:0] \$140 ;
  wire \$142 ;
  wire [8:0] \$144 ;
  wire \$146 ;
  wire [8:0] \$148 ;
  wire \$15 ;
  wire \$150 ;
  wire \$152 ;
  wire \$154 ;
  wire \$156 ;
  wire \$158 ;
  wire \$160 ;
  wire \$162 ;
  wire \$164 ;
  wire \$166 ;
  wire \$168 ;
  wire \$17 ;
  wire \$170 ;
  wire [5:0] \$172 ;
  wire \$174 ;
  wire [5:0] \$176 ;
  wire \$178 ;
  wire [5:0] \$180 ;
  wire \$182 ;
  wire [5:0] \$184 ;
  wire \$186 ;
  wire [5:0] \$188 ;
  wire \$19 ;
  wire \$190 ;
  wire [5:0] \$192 ;
  wire \$194 ;
  wire [5:0] \$196 ;
  wire \$198 ;
  wire [5:0] \$200 ;
  wire \$202 ;
  wire [5:0] \$204 ;
  wire \$206 ;
  wire [5:0] \$208 ;
  wire \$21 ;
  wire \$210 ;
  wire [9:0] \$212 ;
  wire [9:0] \$213 ;
  wire \$215 ;
  wire [5:0] \$217 ;
  wire [6:0] \$219 ;
  wire \$221 ;
  wire [5:0] \$223 ;
  wire [6:0] \$225 ;
  wire \$227 ;
  wire [5:0] \$229 ;
  wire \$23 ;
  wire \$231 ;
  wire \$25 ;
  wire [5:0] \$27 ;
  wire [5:0] \$28 ;
  wire \$3 ;
  wire \$30 ;
  wire [5:0] \$32 ;
  wire [5:0] \$33 ;
  wire \$35 ;
  wire [5:0] \$37 ;
  wire [5:0] \$38 ;
  wire \$40 ;
  wire [5:0] \$42 ;
  wire [5:0] \$43 ;
  wire \$45 ;
  wire [5:0] \$47 ;
  wire [5:0] \$48 ;
  wire \$5 ;
  wire \$50 ;
  wire [5:0] \$52 ;
  wire [5:0] \$53 ;
  wire \$55 ;
  wire [5:0] \$57 ;
  wire [5:0] \$58 ;
  wire \$60 ;
  wire [5:0] \$62 ;
  wire [5:0] \$63 ;
  wire \$65 ;
  wire [5:0] \$67 ;
  wire [5:0] \$68 ;
  wire \$7 ;
  wire \$70 ;
  wire [5:0] \$72 ;
  wire [5:0] \$73 ;
  wire \$75 ;
  wire [5:0] \$77 ;
  wire [5:0] \$78 ;
  wire \$80 ;
  wire [4:0] \$82 ;
  wire [4:0] \$83 ;
  wire \$85 ;
  wire \$87 ;
  wire [3:0] \$89 ;
  wire \$9 ;
  wire [3:0] \$90 ;
  wire [3:0] \$92 ;
  wire [3:0] \$94 ;
  wire [3:0] \$96 ;
  wire [3:0] \$98 ;
  input clk;
  wire clk;
  reg [3:0] curNoteIndex = 4'h0;
  reg [3:0] \curNoteIndex$next ;
  (* enum_base_type = "DiscriminatorState" *)
  (* enum_value_000 = "PowerUp" *)
  (* enum_value_001 = "Init" *)
  (* enum_value_010 = "CalculateDiffFromTarget" *)
  (* enum_value_011 = "Compare" *)
  (* enum_value_100 = "MovedToNextCheckBounds" *)
  (* enum_value_101 = "DetectedValidNote" *)
  (* enum_value_110 = "DisplayResult" *)
  reg [2:0] curState = 3'h0;
  reg [2:0] \curState$next ;
  reg [5:0] detectionWindow = 6'h00;
  reg [5:0] \detectionWindow$next ;
  reg [5:0] detectionWindowMidPoint = 6'h00;
  reg [5:0] \detectionWindowMidPoint$next ;
  input [7:0] edge_count;
  wire [7:0] edge_count;
  reg inputFreqHigher = 1'h0;
  reg \inputFreqHigher$next ;
  output match_exact;
  reg match_exact = 1'h0;
  reg \match_exact$next ;
  output match_far;
  reg match_far = 1'h0;
  reg \match_far$next ;
  output match_high;
  reg match_high = 1'h0;
  reg \match_high$next ;
  reg [4:0] noMatchCount = 5'h00;
  reg [4:0] \noMatchCount$next ;
  output [3:0] note;
  reg [3:0] note = 4'h0;
  reg [3:0] \note$next ;
  reg [5:0] readingProximityResult = 6'h00;
  reg [5:0] \readingProximityResult$next ;
  input rst;
  wire rst;
  reg [8:0] subtractResult = 9'h000;
  reg [8:0] \subtractResult$next ;
  assign \$9  = edge_count > 8'h51;
  assign \$110  = edge_count > 8'h91;
  assign \$112  = 8'h91 - edge_count;
  assign \$114  = edge_count > 8'h7a;
  assign \$116  = 8'h7a - edge_count;
  assign \$118  = edge_count > 8'h6d;
  assign \$11  = edge_count > 8'h49;
  assign \$120  = 8'h6d - edge_count;
  assign \$122  = edge_count > 8'h5b;
  assign \$124  = 8'h5b - edge_count;
  assign \$126  = edge_count > 8'h51;
  assign \$128  = 8'h51 - edge_count;
  assign \$130  = edge_count > 8'h49;
  assign \$132  = 8'h49 - edge_count;
  assign \$134  = edge_count > 8'h3d;
  assign \$136  = 8'h3d - edge_count;
  assign \$138  = edge_count > 8'h36;
  assign \$13  = edge_count > 8'h3d;
  assign \$140  = 8'h36 - edge_count;
  assign \$142  = edge_count > 8'h28;
  assign \$144  = 8'h28 - edge_count;
  assign \$146  = edge_count > 8'h1e;
  assign \$148  = 8'h1e - edge_count;
  assign \$150  = edge_count > 8'h91;
  assign \$152  = edge_count > 8'h7a;
  assign \$154  = edge_count > 8'h6d;
  assign \$156  = edge_count > 8'h5b;
  assign \$158  = edge_count > 8'h51;
  assign \$15  = edge_count > 8'h36;
  assign \$160  = edge_count > 8'h49;
  assign \$162  = edge_count > 8'h3d;
  assign \$164  = edge_count > 8'h36;
  assign \$166  = edge_count > 8'h28;
  assign \$168  = edge_count > 8'h1e;
  assign \$170  = edge_count > 8'h91;
  assign \$174  = edge_count > 8'h7a;
  assign \$178  = edge_count > 8'h6d;
  assign \$17  = edge_count > 8'h28;
  assign \$182  = edge_count > 8'h5b;
  assign \$186  = edge_count > 8'h51;
  assign \$190  = edge_count > 8'h49;
  assign \$194  = edge_count > 8'h3d;
  assign \$198  = edge_count > 8'h36;
  assign \$1  = edge_count > 8'h91;
  assign \$19  = edge_count > 8'h1e;
  assign \$202  = edge_count > 8'h28;
  assign \$206  = edge_count > 8'h1e;
  assign \$210  = subtractResult <= detectionWindowMidPoint;
  assign \$213  = detectionWindow - subtractResult;
  assign \$215  = subtractResult <= detectionWindowMidPoint;
  assign \$21  = subtractResult <= detectionWindow;
  assign \$219  = detectionWindowMidPoint - \$217 ;
  assign \$221  = readingProximityResult >= \$219 ;
  assign \$225  = detectionWindowMidPoint - \$223 ;
  assign \$227  = readingProximityResult >= \$225 ;
  assign \$231  = readingProximityResult <= \$229 ;
  always @(posedge clk)
    curState <= \curState$next ;
  always @(posedge clk)
    noMatchCount <= \noMatchCount$next ;
  always @(posedge clk)
    curNoteIndex <= \curNoteIndex$next ;
  always @(posedge clk)
    note <= \note$next ;
  always @(posedge clk)
    subtractResult <= \subtractResult$next ;
  always @(posedge clk)
    detectionWindow <= \detectionWindow$next ;
  always @(posedge clk)
    detectionWindowMidPoint <= \detectionWindowMidPoint$next ;
  assign \$23  = curNoteIndex < 4'ha;
  always @(posedge clk)
    readingProximityResult <= \readingProximityResult$next ;
  always @(posedge clk)
    inputFreqHigher <= \inputFreqHigher$next ;
  always @(posedge clk)
    match_exact <= \match_exact$next ;
  always @(posedge clk)
    match_far <= \match_far$next ;
  always @(posedge clk)
    match_high <= \match_high$next ;
  assign \$25  = edge_count > 8'h91;
  assign \$28  = noMatchCount + 1'h1;
  assign \$30  = edge_count > 8'h7a;
  assign \$33  = noMatchCount + 1'h1;
  assign \$35  = edge_count > 8'h6d;
  assign \$38  = noMatchCount + 1'h1;
  assign \$3  = edge_count > 8'h7a;
  assign \$40  = edge_count > 8'h5b;
  assign \$43  = noMatchCount + 1'h1;
  assign \$45  = edge_count > 8'h51;
  assign \$48  = noMatchCount + 1'h1;
  assign \$50  = edge_count > 8'h49;
  assign \$53  = noMatchCount + 1'h1;
  assign \$55  = edge_count > 8'h3d;
  assign \$58  = noMatchCount + 1'h1;
  assign \$5  = edge_count > 8'h6d;
  assign \$60  = edge_count > 8'h36;
  assign \$63  = noMatchCount + 1'h1;
  assign \$65  = edge_count > 8'h28;
  assign \$68  = noMatchCount + 1'h1;
  assign \$70  = edge_count > 8'h1e;
  assign \$73  = noMatchCount + 1'h1;
  assign \$75  = curNoteIndex < 4'ha;
  assign \$78  = noMatchCount + 1'h1;
  assign \$7  = edge_count > 8'h5b;
  assign \$80  = subtractResult <= detectionWindow;
  assign \$83  = curNoteIndex + 1'h1;
  assign \$85  = noMatchCount == 5'h1f;
  assign \$87  = subtractResult <= detectionWindow;
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    casez (curState)
      3'h0:
          \curState$next  = 3'h1;
      3'h1:
          \curState$next  = 3'h2;
      3'h2:
          (* full_case = 32'd1 *)
          casez (curNoteIndex)
            4'h0:
                (* full_case = 32'd1 *)
                casez (\$1 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
            4'h1:
                (* full_case = 32'd1 *)
                casez (\$3 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
            4'h2:
                (* full_case = 32'd1 *)
                casez (\$5 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
            4'h3:
                (* full_case = 32'd1 *)
                casez (\$7 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
            4'h4:
                (* full_case = 32'd1 *)
                casez (\$9 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
            4'h5:
                (* full_case = 32'd1 *)
                casez (\$11 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
            4'h6:
                (* full_case = 32'd1 *)
                casez (\$13 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
            4'h7:
                (* full_case = 32'd1 *)
                casez (\$15 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
            4'h8:
                (* full_case = 32'd1 *)
                casez (\$17 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
            4'h?:
                (* full_case = 32'd1 *)
                casez (\$19 )
                  1'h1:
                      \curState$next  = 3'h1;
                  default:
                      \curState$next  = 3'h3;
                endcase
          endcase
      3'h3:
          (* full_case = 32'd1 *)
          casez (\$21 )
            1'h1:
                \curState$next  = 3'h5;
            default:
                \curState$next  = 3'h4;
          endcase
      3'h4:
          (* full_case = 32'd1 *)
          casez (\$23 )
            1'h1:
                \curState$next  = 3'h2;
            default:
                \curState$next  = 3'h1;
          endcase
      3'h5:
          \curState$next  = 3'h6;
      3'h6:
          \curState$next  = 3'h1;
      default:
          \curState$next  = 3'h0;
    endcase
    casez (rst)
      1'h1:
          \curState$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \noMatchCount$next  = noMatchCount;
    casez (curState)
      3'h0:
          \noMatchCount$next  = 5'h00;
      3'h1:
          /* empty */;
      3'h2:
          (* full_case = 32'd1 *)
          casez (curNoteIndex)
            4'h0:
                casez (\$25 )
                  1'h1:
                      \noMatchCount$next  = \$28 [4:0];
                endcase
            4'h1:
                casez (\$30 )
                  1'h1:
                      \noMatchCount$next  = \$33 [4:0];
                endcase
            4'h2:
                casez (\$35 )
                  1'h1:
                      \noMatchCount$next  = \$38 [4:0];
                endcase
            4'h3:
                casez (\$40 )
                  1'h1:
                      \noMatchCount$next  = \$43 [4:0];
                endcase
            4'h4:
                casez (\$45 )
                  1'h1:
                      \noMatchCount$next  = \$48 [4:0];
                endcase
            4'h5:
                casez (\$50 )
                  1'h1:
                      \noMatchCount$next  = \$53 [4:0];
                endcase
            4'h6:
                casez (\$55 )
                  1'h1:
                      \noMatchCount$next  = \$58 [4:0];
                endcase
            4'h7:
                casez (\$60 )
                  1'h1:
                      \noMatchCount$next  = \$63 [4:0];
                endcase
            4'h8:
                casez (\$65 )
                  1'h1:
                      \noMatchCount$next  = \$68 [4:0];
                endcase
            4'h?:
                casez (\$70 )
                  1'h1:
                      \noMatchCount$next  = \$73 [4:0];
                endcase
          endcase
      3'h3:
          /* empty */;
      3'h4:
          (* full_case = 32'd1 *)
          casez (\$75 )
            1'h1:
                /* empty */;
            default:
                \noMatchCount$next  = \$78 [4:0];
          endcase
      3'h5:
          \noMatchCount$next  = 5'h00;
    endcase
    casez (rst)
      1'h1:
          \noMatchCount$next  = 5'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \match_far$next  = match_far;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          /* empty */;
      3'h2:
          /* empty */;
      3'h3:
          /* empty */;
      3'h4:
          /* empty */;
      3'h5:
          /* empty */;
      3'h6:
          (* full_case = 32'd1 *)
          casez (\$227 )
            1'h1:
                \match_far$next  = 1'h0;
            default:
                (* full_case = 32'd1 *)
                casez (\$231 )
                  1'h1:
                      \match_far$next  = 1'h1;
                  default:
                      \match_far$next  = 1'h0;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \match_far$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \match_high$next  = match_high;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          /* empty */;
      3'h2:
          /* empty */;
      3'h3:
          /* empty */;
      3'h4:
          /* empty */;
      3'h5:
          /* empty */;
      3'h6:
          \match_high$next  = inputFreqHigher;
    endcase
    casez (rst)
      1'h1:
          \match_high$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \curNoteIndex$next  = curNoteIndex;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          \curNoteIndex$next  = 4'h0;
      3'h2:
          /* empty */;
      3'h3:
          (* full_case = 32'd1 *)
          casez (\$80 )
            1'h1:
                /* empty */;
            default:
                \curNoteIndex$next  = \$83 [3:0];
          endcase
    endcase
    casez (rst)
      1'h1:
          \curNoteIndex$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \note$next  = note;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          casez (\$85 )
            1'h1:
                \note$next  = 4'h0;
          endcase
      3'h2:
          /* empty */;
      3'h3:
          casez (\$87 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (curNoteIndex)
                  4'h0:
                      \note$next  = \$90 ;
                  4'h1:
                      \note$next  = \$92 ;
                  4'h2:
                      \note$next  = \$94 ;
                  4'h3:
                      \note$next  = \$96 ;
                  4'h4:
                      \note$next  = \$98 ;
                  4'h5:
                      \note$next  = \$100 ;
                  4'h6:
                      \note$next  = \$102 ;
                  4'h7:
                      \note$next  = \$104 ;
                  4'h8:
                      \note$next  = \$106 ;
                  4'h?:
                      \note$next  = \$108 ;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \note$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \subtractResult$next  = subtractResult;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          /* empty */;
      3'h2:
          (* full_case = 32'd1 *)
          casez (curNoteIndex)
            4'h0:
                (* full_case = 32'd1 *)
                casez (\$110 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$112 ;
                endcase
            4'h1:
                (* full_case = 32'd1 *)
                casez (\$114 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$116 ;
                endcase
            4'h2:
                (* full_case = 32'd1 *)
                casez (\$118 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$120 ;
                endcase
            4'h3:
                (* full_case = 32'd1 *)
                casez (\$122 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$124 ;
                endcase
            4'h4:
                (* full_case = 32'd1 *)
                casez (\$126 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$128 ;
                endcase
            4'h5:
                (* full_case = 32'd1 *)
                casez (\$130 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$132 ;
                endcase
            4'h6:
                (* full_case = 32'd1 *)
                casez (\$134 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$136 ;
                endcase
            4'h7:
                (* full_case = 32'd1 *)
                casez (\$138 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$140 ;
                endcase
            4'h8:
                (* full_case = 32'd1 *)
                casez (\$142 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$144 ;
                endcase
            4'h?:
                (* full_case = 32'd1 *)
                casez (\$146 )
                  1'h1:
                      /* empty */;
                  default:
                      \subtractResult$next  = \$148 ;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \subtractResult$next  = 9'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \detectionWindow$next  = detectionWindow;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          /* empty */;
      3'h2:
          (* full_case = 32'd1 *)
          casez (curNoteIndex)
            4'h0:
                (* full_case = 32'd1 *)
                casez (\$150 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h11;
                endcase
            4'h1:
                (* full_case = 32'd1 *)
                casez (\$152 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h0e;
                endcase
            4'h2:
                (* full_case = 32'd1 *)
                casez (\$154 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h0c;
                endcase
            4'h3:
                (* full_case = 32'd1 *)
                casez (\$156 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h0a;
                endcase
            4'h4:
                (* full_case = 32'd1 *)
                casez (\$158 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h09;
                endcase
            4'h5:
                (* full_case = 32'd1 *)
                casez (\$160 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h08;
                endcase
            4'h6:
                (* full_case = 32'd1 *)
                casez (\$162 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h07;
                endcase
            4'h7:
                (* full_case = 32'd1 *)
                casez (\$164 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h06;
                endcase
            4'h8:
                (* full_case = 32'd1 *)
                casez (\$166 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h04;
                endcase
            4'h?:
                (* full_case = 32'd1 *)
                casez (\$168 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindow$next  = 6'h03;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \detectionWindow$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \detectionWindowMidPoint$next  = detectionWindowMidPoint;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          /* empty */;
      3'h2:
          (* full_case = 32'd1 *)
          casez (curNoteIndex)
            4'h0:
                (* full_case = 32'd1 *)
                casez (\$170 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$172 ;
                endcase
            4'h1:
                (* full_case = 32'd1 *)
                casez (\$174 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$176 ;
                endcase
            4'h2:
                (* full_case = 32'd1 *)
                casez (\$178 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$180 ;
                endcase
            4'h3:
                (* full_case = 32'd1 *)
                casez (\$182 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$184 ;
                endcase
            4'h4:
                (* full_case = 32'd1 *)
                casez (\$186 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$188 ;
                endcase
            4'h5:
                (* full_case = 32'd1 *)
                casez (\$190 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$192 ;
                endcase
            4'h6:
                (* full_case = 32'd1 *)
                casez (\$194 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$196 ;
                endcase
            4'h7:
                (* full_case = 32'd1 *)
                casez (\$198 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$200 ;
                endcase
            4'h8:
                (* full_case = 32'd1 *)
                casez (\$202 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$204 ;
                endcase
            4'h?:
                (* full_case = 32'd1 *)
                casez (\$206 )
                  1'h1:
                      /* empty */;
                  default:
                      \detectionWindowMidPoint$next  = \$208 ;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \detectionWindowMidPoint$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \readingProximityResult$next  = readingProximityResult;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          /* empty */;
      3'h2:
          /* empty */;
      3'h3:
          /* empty */;
      3'h4:
          /* empty */;
      3'h5:
          (* full_case = 32'd1 *)
          casez (\$210 )
            1'h1:
                \readingProximityResult$next  = subtractResult[5:0];
            default:
                \readingProximityResult$next  = \$213 [5:0];
          endcase
    endcase
    casez (rst)
      1'h1:
          \readingProximityResult$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \inputFreqHigher$next  = inputFreqHigher;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          /* empty */;
      3'h2:
          /* empty */;
      3'h3:
          /* empty */;
      3'h4:
          /* empty */;
      3'h5:
          (* full_case = 32'd1 *)
          casez (\$215 )
            1'h1:
                \inputFreqHigher$next  = 1'h1;
            default:
                \inputFreqHigher$next  = 1'h0;
          endcase
    endcase
    casez (rst)
      1'h1:
          \inputFreqHigher$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$5 ) begin end
    \match_exact$next  = match_exact;
    casez (curState)
      3'h0:
          /* empty */;
      3'h1:
          /* empty */;
      3'h2:
          /* empty */;
      3'h3:
          /* empty */;
      3'h4:
          /* empty */;
      3'h5:
          /* empty */;
      3'h6:
          (* full_case = 32'd1 *)
          casez (\$221 )
            1'h1:
                \match_exact$next  = 1'h1;
            default:
                \match_exact$next  = 1'h0;
          endcase
    endcase
    casez (rst)
      1'h1:
          \match_exact$next  = 1'h0;
    endcase
  end
  assign \$27  = \$28 ;
  assign \$32  = \$33 ;
  assign \$37  = \$38 ;
  assign \$42  = \$43 ;
  assign \$47  = \$48 ;
  assign \$52  = \$53 ;
  assign \$57  = \$58 ;
  assign \$62  = \$63 ;
  assign \$67  = \$68 ;
  assign \$72  = \$73 ;
  assign \$77  = \$78 ;
  assign \$82  = \$83 ;
  assign \$212  = \$213 ;
  assign \$90  = 4'h1;
  assign \$92  = 4'h6;
  assign \$94  = 4'h5;
  assign \$96  = 4'h3;
  assign \$98  = 4'h2;
  assign \$100  = 4'h1;
  assign \$102  = 4'h6;
  assign \$104  = 4'h5;
  assign \$106  = 4'h2;
  assign \$108  = 4'h6;
  assign \$172  = 6'h08;
  assign \$176  = 6'h07;
  assign \$180  = 6'h06;
  assign \$184  = 6'h05;
  assign \$188  = 6'h04;
  assign \$192  = 6'h04;
  assign \$196  = 6'h03;
  assign \$200  = 6'h03;
  assign \$204  = 6'h02;
  assign \$208  = 6'h01;
  assign \$217  = { 4'h0, detectionWindow[5:4] };
  assign \$223  = { 4'h0, detectionWindow[5:4] };
  assign \$229  = { 1'h0, detectionWindowMidPoint[5:1] };
endmodule

module display(clk, valueNote, valueProxim, segments, proximitySelect, rst);
  reg \$auto$verilog_backend.cc:2097:dump_module$6  = 0;
  wire \$1 ;
  input clk;
  wire clk;
  wire [7:0] notedisplay_segments;
  reg [2:0] notedisplay_value = 3'h0;
  reg [2:0] \notedisplay_value$next ;
  wire [7:0] proxdisplay_segments;
  reg [2:0] proxdisplay_value = 3'h0;
  reg [2:0] \proxdisplay_value$next ;
  output proximitySelect;
  reg proximitySelect = 1'h0;
  reg \proximitySelect$next ;
  input rst;
  wire rst;
  output [7:0] segments;
  reg [7:0] segments = 8'h00;
  reg [7:0] \segments$next ;
  input [3:0] valueNote;
  wire [3:0] valueNote;
  input [2:0] valueProxim;
  wire [2:0] valueProxim;
  assign \$1  = ! valueNote;
  always @(posedge clk)
    notedisplay_value <= \notedisplay_value$next ;
  always @(posedge clk)
    proxdisplay_value <= \proxdisplay_value$next ;
  always @(posedge clk)
    proximitySelect <= \proximitySelect$next ;
  always @(posedge clk)
    segments <= \segments$next ;
  notedisplay notedisplay (
    .clk(clk),
    .rst(rst),
    .segments(notedisplay_segments),
    .value(notedisplay_value)
  );
  proxdisplay proxdisplay (
    .clk(clk),
    .rst(rst),
    .segments(proxdisplay_segments),
    .value(proxdisplay_value)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$6 ) begin end
    \notedisplay_value$next  = valueNote[2:0];
    casez (rst)
      1'h1:
          \notedisplay_value$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$6 ) begin end
    \proxdisplay_value$next  = valueProxim;
    casez (rst)
      1'h1:
          \proxdisplay_value$next  = 3'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$6 ) begin end
    \proximitySelect$next  = 1'h1;
    casez (proximitySelect)
      1'h1:
          \proximitySelect$next  = 1'h0;
    endcase
    casez (rst)
      1'h1:
          \proximitySelect$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$6 ) begin end
    (* full_case = 32'd1 *)
    casez (proximitySelect)
      1'h1:
          (* full_case = 32'd1 *)
          casez (\$1 )
            1'h1:
                \segments$next  = notedisplay_segments;
            default:
                \segments$next  = proxdisplay_segments;
          endcase
      default:
          \segments$next  = notedisplay_segments;
    endcase
    casez (rst)
      1'h1:
          \segments$next  = 8'h00;
    endcase
  end
endmodule

module edge_detect(clk, \input , \output , rst);
  reg \$auto$verilog_backend.cc:2097:dump_module$7  = 0;
  wire \$1 ;
  wire \$3 ;
  input clk;
  wire clk;
  wire ffsync_syncOut;
  input \input ;
  wire \input ;
  output \output ;
  reg \output  = 1'h0;
  reg \output$next ;
  input rst;
  wire rst;
  reg seenRising = 1'h0;
  reg \seenRising$next ;
  assign \$1  = ~ seenRising;
  assign \$3  = ~ seenRising;
  always @(posedge clk)
    \output  <= \output$next ;
  always @(posedge clk)
    seenRising <= \seenRising$next ;
  ffsync ffsync (
    .clk(clk),
    .\input (\input ),
    .rst(rst),
    .syncOut(ffsync_syncOut)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$7 ) begin end
    \output$next  = 1'h0;
    casez (ffsync_syncOut)
      1'h1:
          casez (\$1 )
            1'h1:
                \output$next  = 1'h1;
          endcase
    endcase
    casez (rst)
      1'h1:
          \output$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$7 ) begin end
    \seenRising$next  = seenRising;
    (* full_case = 32'd1 *)
    casez (ffsync_syncOut)
      1'h1:
          casez (\$3 )
            1'h1:
                \seenRising$next  = 1'h1;
          endcase
      default:
          \seenRising$next  = 1'h0;
    endcase
    casez (rst)
      1'h1:
          \seenRising$next  = 1'h0;
    endcase
  end
endmodule

module ffsync(clk, \input , syncOut, rst);
  input clk;
  wire clk;
  input \input ;
  wire \input ;
  input rst;
  wire rst;
  reg stage0 = 1'h0;
  wire \stage0$next ;
  reg stage1 = 1'h0;
  wire \stage1$next ;
  output syncOut;
  wire syncOut;
  always @(posedge clk)
    stage0 <= \stage0$next ;
  always @(posedge clk)
    stage1 <= \stage1$next ;
  assign syncOut = stage1;
  assign \stage1$next  = stage0;
  assign \stage0$next  = \input ;
endmodule

module notedisplay(clk, value, segments, rst);
  reg \$auto$verilog_backend.cc:2097:dump_module$8  = 0;
  wire \$1 ;
  input clk;
  wire clk;
  input rst;
  wire rst;
  output [7:0] segments;
  reg [7:0] segments = 8'h00;
  reg [7:0] \segments$next ;
  input [2:0] value;
  wire [2:0] value;
  assign \$1  = value < 4'h8;
  always @(posedge clk)
    segments <= \segments$next ;
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$8 ) begin end
    \segments$next  = 8'h00;
    casez (\$1 )
      1'h1:
          (* full_case = 32'd1 *)
          casez (value)
            3'h0:
                \segments$next  = 8'h02;
            3'h1:
                \segments$next  = 8'hf6;
            3'h2:
                \segments$next  = 8'hee;
            3'h3:
                \segments$next  = 8'h3e;
            3'h4:
                \segments$next  = 8'h9c;
            3'h5:
                \segments$next  = 8'h7a;
            3'h6:
                \segments$next  = 8'h9e;
            3'h?:
                \segments$next  = 8'h8e;
          endcase
    endcase
    casez (rst)
      1'h1:
          \segments$next  = 8'h00;
    endcase
  end
endmodule

module proxdisplay(clk, value, segments, rst);
  reg \$auto$verilog_backend.cc:2097:dump_module$9  = 0;
  wire \$1 ;
  input clk;
  wire clk;
  input rst;
  wire rst;
  output [7:0] segments;
  reg [7:0] segments = 8'h00;
  reg [7:0] \segments$next ;
  input [2:0] value;
  wire [2:0] value;
  assign \$1  = value < 4'h8;
  always @(posedge clk)
    segments <= \segments$next ;
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$9 ) begin end
    \segments$next  = 8'h00;
    casez (\$1 )
      1'h1:
          (* full_case = 32'd1 *)
          casez (value)
            3'h0:
                \segments$next  = 8'h2a;
            3'h1:
                \segments$next  = 8'h01;
            3'h2:
                \segments$next  = 8'h46;
            3'h3:
                \segments$next  = 8'h01;
            3'h4:
                \segments$next  = 8'h38;
            3'h5:
                \segments$next  = 8'h01;
            3'h6:
                \segments$next  = 8'hc4;
            3'h?:
                \segments$next  = 8'h01;
          endcase
    endcase
    casez (rst)
      1'h1:
          \segments$next  = 8'h00;
    endcase
  end
endmodule

module pulsecounter(clk, \input , clock_config, pulseCount, rst);
  reg \$auto$verilog_backend.cc:2097:dump_module$10  = 0;
  wire [15:0] \$1 ;
  wire \$10 ;
  wire [15:0] \$12 ;
  wire [15:0] \$13 ;
  wire [15:0] \$2 ;
  wire \$4 ;
  wire \$6 ;
  wire \$8 ;
  wire [14:0] \$auto$proc_rom.cc:149:do_switch$1 ;
  input clk;
  wire clk;
  reg [14:0] clockCount = 15'h0000;
  reg [14:0] \clockCount$next ;
  input [2:0] clock_config;
  wire [2:0] clock_config;
  wire edge_detect_input;
  wire edge_detect_output;
  input \input ;
  wire \input ;
  output [14:0] pulseCount;
  reg [14:0] pulseCount = 15'h0000;
  reg [14:0] \pulseCount$next ;
  input rst;
  wire rst;
  reg [14:0] runningPulseCount = 15'h0000;
  reg [14:0] \runningPulseCount$next ;
  reg [14:0] singlePeriodClockCount = 15'h0000;
  reg [14:0] \singlePeriodClockCount$next ;
  (* full_case = 32'd1 *)
  reg [14:0] \$auto$proc_rom.cc:150:do_switch$2  [7:0];
  initial begin
    \$auto$proc_rom.cc:150:do_switch$2 [0] = 15'h015e;
    \$auto$proc_rom.cc:150:do_switch$2 [1] = 15'h02bc;
    \$auto$proc_rom.cc:150:do_switch$2 [2] = 15'h0578;
    \$auto$proc_rom.cc:150:do_switch$2 [3] = 15'h047b;
    \$auto$proc_rom.cc:150:do_switch$2 [4] = 15'h0dac;
    \$auto$proc_rom.cc:150:do_switch$2 [5] = 15'h2ccd;
    \$auto$proc_rom.cc:150:do_switch$2 [6] = 15'h36b0;
    \$auto$proc_rom.cc:150:do_switch$2 [7] = 15'h5208;
  end
  assign \$auto$proc_rom.cc:149:do_switch$1  = \$auto$proc_rom.cc:150:do_switch$2 [clock_config];
  assign \$10  = ! clockCount;
  assign \$13  = runningPulseCount + 1'h1;
  always @(posedge clk)
    clockCount <= \clockCount$next ;
  always @(posedge clk)
    singlePeriodClockCount <= \singlePeriodClockCount$next ;
  always @(posedge clk)
    pulseCount <= \pulseCount$next ;
  always @(posedge clk)
    runningPulseCount <= \runningPulseCount$next ;
  assign \$2  = clockCount + 1'h1;
  assign \$4  = clockCount == singlePeriodClockCount;
  assign \$6  = clockCount == singlePeriodClockCount;
  assign \$8  = clockCount == singlePeriodClockCount;
  edge_detect edge_detect (
    .clk(clk),
    .\input (edge_detect_input),
    .\output (edge_detect_output),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$10 ) begin end
    \clockCount$next  = \$2 [14:0];
    casez (\$4 )
      1'h1:
          \clockCount$next  = 15'h0000;
    endcase
    casez (rst)
      1'h1:
          \clockCount$next  = 15'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$10 ) begin end
    \singlePeriodClockCount$next  = \$auto$proc_rom.cc:149:do_switch$1 ;
    casez (rst)
      1'h1:
          \singlePeriodClockCount$next  = 15'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$10 ) begin end
    \pulseCount$next  = pulseCount;
    casez (\$6 )
      1'h1:
          \pulseCount$next  = runningPulseCount;
    endcase
    casez (rst)
      1'h1:
          \pulseCount$next  = 15'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$10 ) begin end
    \runningPulseCount$next  = runningPulseCount;
    (* full_case = 32'd1 *)
    casez (\$8 )
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$10 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (edge_detect_output)
                  1'h1:
                      \runningPulseCount$next  = 15'h0001;
                  default:
                      \runningPulseCount$next  = 15'h0000;
                endcase
            default:
                casez (edge_detect_output)
                  1'h1:
                      \runningPulseCount$next  = \$13 [14:0];
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \runningPulseCount$next  = 15'h0000;
    endcase
  end
  assign \$1  = \$2 ;
  assign \$12  = \$13 ;
  assign edge_detect_input = \input ;
endmodule

module tt_um_psychogenic_neptuneproportional(uo_out, uio_in, uio_out, uio_oe, ena, clk, rst_n, \clk$1 , rst, ui_in);
  reg \$auto$verilog_backend.cc:2097:dump_module$11  = 0;
  input clk;
  wire clk;
  input \clk$1 ;
  wire \clk$1 ;
  reg [7:0] displaySegmentsA = 8'h00;
  reg [7:0] \displaySegmentsA$next ;
  reg [7:0] displaySegmentsB = 8'h00;
  reg [7:0] \displaySegmentsB$next ;
  input ena;
  wire ena;
  wire input_pulses;
  reg [7:0] outputs;
  input rst;
  wire rst;
  input rst_n;
  wire rst_n;
  wire [2:0] tuner_clock_config;
  wire [7:0] tuner_displaySegments;
  wire tuner_displaySelect;
  wire tuner_input_pulses;
  wire tuner_match_exact;
  wire [7:0] tuner_pulseCount;
  input [7:0] ui_in;
  wire [7:0] ui_in;
  input [7:0] uio_in;
  wire [7:0] uio_in;
  output [7:0] uio_oe;
  wire [7:0] uio_oe;
  output [7:0] uio_out;
  wire [7:0] uio_out;
  output [7:0] uo_out;
  wire [7:0] uo_out;
  always @(posedge \clk$1 )
    displaySegmentsA <= \displaySegmentsA$next ;
  always @(posedge \clk$1 )
    displaySegmentsB <= \displaySegmentsB$next ;
  tuner tuner (
    .clk(\clk$1 ),
    .clock_config(tuner_clock_config),
    .displaySegments(tuner_displaySegments),
    .displaySelect(tuner_displaySelect),
    .input_pulses(tuner_input_pulses),
    .match_exact(tuner_match_exact),
    .pulseCount(tuner_pulseCount),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$11 ) begin end
    \displaySegmentsA$next  = displaySegmentsA;
    casez (tuner_displaySelect)
      1'h1:
          \displaySegmentsA$next  = { tuner_displaySegments[7:1], tuner_match_exact };
    endcase
    casez (rst)
      1'h1:
          \displaySegmentsA$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$11 ) begin end
    \displaySegmentsB$next  = displaySegmentsB;
    (* full_case = 32'd1 *)
    casez (tuner_displaySelect)
      1'h1:
          /* empty */;
      default:
          \displaySegmentsB$next  = tuner_displaySegments;
    endcase
    casez (rst)
      1'h1:
          \displaySegmentsB$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$11 ) begin end
    (* full_case = 32'd1 *)
    casez (ui_in[6])
      1'h1:
          (* full_case = 32'd1 *)
          casez (ui_in[7])
            1'h1:
                outputs = displaySegmentsA;
            default:
                outputs = displaySegmentsB;
          endcase
      default:
          outputs = { tuner_displaySelect, tuner_displaySegments[7:1] };
    endcase
  end
  assign uo_out = outputs;
  assign tuner_input_pulses = ui_in[5];
  assign tuner_clock_config = ui_in[4:2];
  assign input_pulses = ui_in[5];
  assign uio_out = tuner_pulseCount;
  assign uio_oe = 8'hff;
endmodule

module tuner(clock_config, input_pulses, displaySelect, match_exact, displaySegments, rst, clk, pulseCount);
  input clk;
  wire clk;
  input [2:0] clock_config;
  wire [2:0] clock_config;
  wire [7:0] discriminator_edge_count;
  wire discriminator_match_far;
  wire discriminator_match_high;
  wire [3:0] discriminator_note;
  output [7:0] displaySegments;
  wire [7:0] displaySegments;
  output displaySelect;
  wire displaySelect;
  wire display_proximitySelect;
  wire [7:0] display_segments;
  wire [3:0] display_valueNote;
  wire [2:0] display_valueProxim;
  input input_pulses;
  wire input_pulses;
  output match_exact;
  wire match_exact;
  output [7:0] pulseCount;
  wire [7:0] pulseCount;
  wire [2:0] pulsecounter_clock_config;
  wire pulsecounter_input;
  wire [14:0] pulsecounter_pulseCount;
  input rst;
  wire rst;
  discriminator discriminator (
    .clk(clk),
    .edge_count(discriminator_edge_count),
    .match_exact(match_exact),
    .match_far(discriminator_match_far),
    .match_high(discriminator_match_high),
    .note(discriminator_note),
    .rst(rst)
  );
  display display (
    .clk(clk),
    .proximitySelect(display_proximitySelect),
    .rst(rst),
    .segments(display_segments),
    .valueNote(display_valueNote),
    .valueProxim(display_valueProxim)
  );
  pulsecounter pulsecounter (
    .clk(clk),
    .clock_config(pulsecounter_clock_config),
    .\input (pulsecounter_input),
    .pulseCount(pulsecounter_pulseCount),
    .rst(rst)
  );
  assign pulseCount = pulsecounter_pulseCount[7:0];
  assign displaySelect = display_proximitySelect;
  assign displaySegments = display_segments;
  assign display_valueProxim = { discriminator_match_far, discriminator_match_high, match_exact };
  assign display_valueNote = discriminator_note;
  assign discriminator_edge_count = pulsecounter_pulseCount[7:0];
  assign pulsecounter_clock_config = clock_config;
  assign pulsecounter_input = input_pulses;
endmodule

